library verilog;
use verilog.vl_types.all;
entity testAlu is
end testAlu;
