library verilog;
use verilog.vl_types.all;
entity fsm is
    port(
        IR              : in     vl_logic_vector(31 downto 0);
        stat            : out    vl_logic_vector(3 downto 0)
    );
end fsm;
