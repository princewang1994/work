library verilog;
use verilog.vl_types.all;
entity testCtr is
end testCtr;
