library verilog;
use verilog.vl_types.all;
entity testDm is
end testDm;
