library verilog;
use verilog.vl_types.all;
entity test_mul is
end test_mul;
