library verilog;
use verilog.vl_types.all;
entity mux is
end mux;
