library verilog;
use verilog.vl_types.all;
entity mips55 is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end mips55;
