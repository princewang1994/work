library verilog;
use verilog.vl_types.all;
entity testIm is
end testIm;
