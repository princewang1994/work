library verilog;
use verilog.vl_types.all;
entity testext is
end testext;
