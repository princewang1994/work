module cp0(A1,A2,A3,WD1,WD2,CP0Wr,clk,reset,RD);
  
  input [4:0] A1;
  input [4:0] A2;
  input [4:0] A3;
  
  input [31:0]WD1;
  
  input [31:0]WD2;
  
  input [1:0] CP0Wr;
  
  input reset;
  
  input clk;
  
  output [31:0] RD;
  
  reg [31:0] RF[31:0];//reg file;
  
  assign RD=RF[A1];
  
  integer i;
  
  always@(posedge clk)
  begin
    if(reset)
    begin
          for(i=0;i<=31;i=i+1) 
            RF[i]<=0; 
    end
    
    else
    begin
      if(CP0Wr[1])
        RF[A2] <= WD1; 
      if(CP0Wr[0])     
        RF[A3] <= WD2;
    end 

  end
  
  initial
  begin
        for(i=0;i<=31;i=i+1) 
            RF[i]<=0; 
  end
  
  
endmodule


