library verilog;
use verilog.vl_types.all;
entity testmux is
end testmux;
